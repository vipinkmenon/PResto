module or_gate(
input [5:0] I2,
output O2
);

assign O2 = |I2;

endmodule

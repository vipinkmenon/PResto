module and_gate(
input [5:0] I1,
output O1
);

assign O1 = &I1;

endmodule
